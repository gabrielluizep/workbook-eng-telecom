pll5khz_inst : pll5khz PORT MAP (
		inclk0	 => inclk0_sig,
		c0	 => c0_sig
	);
